library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library pll;
use pll.all;

entity telecran is
    port (
        -- FPGA
        i_clk_50: in std_logic;

        -- HDMI
        io_hdmi_i2c_scl       : inout std_logic;
        io_hdmi_i2c_sda       : inout std_logic;
        o_hdmi_tx_clk        : out std_logic;
        o_hdmi_tx_d          : out std_logic_vector(23 downto 0);
        o_hdmi_tx_de         : out std_logic;
        o_hdmi_tx_hs         : out std_logic;
        i_hdmi_tx_int        : in std_logic;
        o_hdmi_tx_vs         : out std_logic;

        -- KEYs
        i_rst_n : in std_logic;
		  
		-- LEDs
		o_leds : out std_logic_vector(9 downto 0);
		o_de10_leds : out std_logic_vector(7 downto 0);

		-- Coder
		i_left_ch_a : in std_logic;
		i_left_ch_b : in std_logic;
		i_left_pb : in std_logic;
		i_right_ch_a : in std_logic;
		i_right_ch_b : in std_logic;
		i_right_pb : in std_logic
    );
end entity telecran;

architecture rtl of telecran is
	component I2C_HDMI_Config 
		port (
			iCLK : in std_logic;
			iRST_N : in std_logic;
			I2C_SCLK : out std_logic;
			I2C_SDAT : inout std_logic;
			HDMI_TX_INT  : in std_logic
		);
	 end component;
	 
	component pll 
		port (
			refclk : in std_logic;
			rst : in std_logic;
			outclk_0 : out std_logic;
			locked : out std_logic
		);
	end component;

    constant h_res : natural := 720;
    constant v_res : natural := 480;
	 

	signal s_clk_27 : std_logic;
	signal s_rst_n : std_logic;	-- holds reset as long as pll is not locked
	
	signal s_x_counter : natural range 0 to h_res - 1;
   signal s_y_counter : natural range 0 to v_res - 1;
	
	signal s_x_encoder : natural range 0 to h_res-1 := 0;
   signal s_y_encoder : natural range 0 to v_res-1 := 0;
	
	signal s_pixel_addr_a : natural range 0 to h_res*v_res-1;
	signal s_pixel_addr_b : natural range 0 to h_res*v_res-1;
	
	signal s_data_a : std_logic_vector(8-1 downto 0);
	signal s_data_out : std_logic_vector(8-1 downto 0);
	
	signal s_clear_flag : std_logic := '0';
	signal s_clear_addr : natural range 0 to h_res*v_res-1 := 0;

begin
	-- o_leds <= (others => '0');
	-- o_de10_leds <= (others => '0');
	
	-- Frequency for HDMI is 27MHz generated by this PLL
	pll0 : component pll 
		port map (
			refclk => i_clk_50,
			rst => not(i_rst_n),
			outclk_0 => s_clk_27,
			locked => s_rst_n
		);

	-- Configures the ADV7513 for 480p
	I2C_HDMI_Config0 : component I2C_HDMI_Config 
		port map (
			iCLK => i_clk_50,
			iRST_N => i_rst_n,
			I2C_SCLK => io_hdmi_i2c_scl,
			I2C_SDAT => io_hdmi_i2c_sda,
			HDMI_TX_INT => i_hdmi_tx_int
	 );
	 
	encodeur_left : entity work.encodeur
	   generic map (
			CNT_MAX => h_res
		)
		port map (
			i_clk => i_clk_50,
			i_rst_n => i_rst_n,
			i_ch_a => i_left_ch_a,
			i_ch_b => i_left_ch_b,
			i_pb => i_left_pb,
			
			o_compteur => s_x_encoder
	);
	
	encodeur_right : entity work.encodeur
		generic map (
			CNT_MAX => v_res
		)
		port map (
			i_clk => i_clk_50,
			i_rst_n => i_rst_n,
			i_ch_a => i_right_ch_a,
			i_ch_b => i_right_ch_b,
			i_pb => i_right_pb,
			
			o_compteur => s_y_encoder
	);
	
	hdmi_controler0 : entity work.hdmi_controler
		port map (
			i_clk => s_clk_27,
			i_rst_n => s_rst_n,
			
			o_hdmi_hs => o_hdmi_tx_hs,
			o_hdmi_vs => o_hdmi_tx_vs,
			o_hdmi_de => o_hdmi_tx_de,
			
			o_pixel_en => open,
			o_pixel_address => s_pixel_addr_b,
			o_x_counter => s_x_counter,
         o_y_counter => s_y_counter
			
	);
	
	dpram0 : entity work.dpram
		generic map (
			mem_size => h_res * v_res,
			data_width => 8
		)
		port map (
		  i_clk_a => i_clk_50,
        i_clk_b => s_clk_27,

        i_data_a => s_data_a,
        i_data_b => x"00",
        i_addr_a => s_pixel_addr_a,
        i_addr_b => s_pixel_addr_b,
        i_we_a => '1',
        i_we_b => '0',
        o_q_a => open,
        o_q_b => s_data_out
	);
	
	o_hdmi_tx_clk <= s_clk_27;
	

	process(i_clk_50)
	begin 
		if rising_edge(i_clk_50) then
		
			if (i_right_pb = '0') then
				s_clear_flag <= '1';
				s_clear_addr <= 0;
				
			end if; 
			
			if (s_clear_flag = '1') then 
				s_pixel_addr_a <= s_clear_addr;
				s_data_a <= x"00";
				
				if (s_clear_addr = h_res*v_res-1) then 
					s_clear_flag <= '0';
					s_clear_addr <= 0;
				else 
					s_clear_addr <= s_clear_addr + 1;
				
				end if;
			else 
				s_pixel_addr_a <= s_x_encoder + (s_y_encoder * h_res);
				s_data_a <= x"FF";
				
			end if;
		end if;
		
	
	end process;
	
	o_hdmi_tx_d(23 downto 16) <= s_data_out;
	
	
end architecture rtl;
